module CLKGT_9T1X ( CK, E, Z);
input  CK;
input  E;
output Z;



endmodule



